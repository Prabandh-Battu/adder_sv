class monitor;
  
  virtual intf vif;
  
  mailbox mon2scb;
  
  function new (virtual intf vif, mailbox mon2scb);
    
    this.vif = vif;
    
    this.mon2scb = mon2scb;
    
  endfunction
  
  task main;
    
    forever begin
      
      transaction trans;
      
      trans = new();
      
      @(posedge vif.clk);
      
      wait(vif.valid);
      
      trans.a <= vif.a;
      
      trans.b <= vif.b;
      
      @(posedge vif.clk);
      
      trans.c = vif.c;
      
      @(posedge vif.clk);
      
      mon2scb.put(trans);
      
      trans.display(":::[MONITOR]:::");
      
    end
    
  endtask
  
endclass
      
      